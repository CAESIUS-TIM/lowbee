`include "../util/util.v"
module test (a);
output a;
reg [util.get_width(5):0] a;    

endmodule