module uart (
    ports
);
    
endmodule